module not_gate(a,y);

input a;
output y;

mux mux1(1'b1,1'b0,a,y);


endmodule

`include "sync_reset.v"
`include "tx.sv"
`include "common.sv"
`include "intf.sv"
`include "gen.sv"
`include "bfm.sv"
`include "agent.sv"
`include "env.sv"
`include "top.sv"
